module inv_22(

	input wire signed [23:0] a,b,c,d,

	output reg signed [23:0] b11,b12,b21,b22
);

reg [23:0] w=24'b0000_0000_1000_0000_0000_0000;
reg signed [47:0] q1,q2,q3,q4;
reg signed [23:0] w1,w2,w3;
reg signed [39:0] w4;

always @(*) 
begin
    w4=w<<15;
    q1=a*d;
    q2={{16{q1[47]}},q1[46:14]};
    q3=b*c;
    q4={{16{q3[47]}},q3[46:14]};
    w1=q2[23:0];
    w2=q4[23:0];
    w3=w1-w2;
    w1=w4/w3; 
    q1=d*w1;
    q2={{16{q1[47]}},q1[46:14]};
    b11=q2[23:0];
    
    q1=a*d;
    q2={{16{q1[47]}},q1[46:14]};
    q3=b*c;
    q4={{16{q3[47]}},q3[46:14]};
    w1=q2[23:0];
    w2=q4[23:0];
    w3=w2-w1;
    w1=w4/w3; 
    q1=b*w1;
    q2={{16{q1[47]}},q1[46:14]};
    b12=q2[23:0];
    
    q1=a*d;
    q2={{16{q1[47]}},q1[46:14]};
    q3=b*c;
    q4={{16{q3[47]}},q3[46:14]};
    w1=q2[23:0];
    w2=q4[23:0];
    w3=w2-w1;
    w1=w4/w3; 
    q1=c*w1;
    q2={{16{q1[47]}},q1[46:14]};
    b21=q2[23:0];
    
    q1=a*d;
    q2={{16{q1[47]}},q1[46:14]};
    q3=b*c;
    q4={{16{q3[47]}},q3[46:14]};
    w1=q2[23:0];
    w2=q4[23:0];
    w3=w1-w2;
    w1=w4/w3; 
    q1=a*w1;
    q2={{16{q1[47]}},q1[46:14]};
    b22=q2[23:0];

end
endmodule
