
module ml_44(
	input wire clk,rst_n,
	input wire signed [23:0] a11,a12,a13,a14,a21,a22,a23,a24,a31,a32,a33,a34,a41,a42,a43,a44,
	input wire signed [23:0] b11,b12,b13,b14,b21,b22,b23,b24,b31,b32,b33,b34,b41,b42,b43,b44,
	output reg signed [23:0] c11,c12,c13,c14,c21,c22,c23,c24,c31,c32,c33,c34,c41,c42,c43,c44 
);

reg signed [47:0] q1,q2,q3,q4,q5;
reg signed [23:0] w1,w2,w3,w4;

always @(clk or ~rst_n ) 
begin
    q1=a11*b11;
    q2=a12*b21;
    q3=a13*b31;
    q4=a14*b41;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c11=w1+w2+w3+w4;
    
    q1=a11*b12;
    q2=a12*b22;
    q3=a13*b32;
    q4=a14*b42;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c12=w1+w2+w3+w4;
    
    q1=a11*b13;
    q2=a12*b23;
    q3=a13*b33;
    q4=a14*b43;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c13=w1+w2+w3+w4;
    
    q1=a11*b14;
    q2=a12*b24;
    q3=a13*b34;
    q4=a14*b44;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c14=w1+w2+w3+w4;
    
    q1=a21*b11;
    q2=a22*b21;
    q3=a23*b31;
    q4=a24*b41;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c21=w1+w2+w3+w4;
    
    q1=a21*b12;
    q2=a22*b22;
    q3=a23*b32;
    q4=a24*b42;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c22=w1+w2+w3+w4;
    
    q1=a21*b13;
    q2=a22*b23;
    q3=a23*b33;
    q4=a24*b43;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c23=w1+w2+w3+w4;
    
    q1=a21*b14;
    q2=a22*b24;
    q3=a23*b34;
    q4=a24*b44;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c24=w1+w2+w3+w4;
    
    q1=a31*b11;
    q2=a32*b21;
    q3=a33*b31;
    q4=a34*b41;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c31=w1+w2+w3+w4;
    
    q1=a31*b12;
    q2=a32*b22;
    q3=a33*b32;
    q4=a34*b42;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c32=w1+w2+w3+w4;
    
    q1=a31*b13;
    q2=a32*b23;
    q3=a33*b33;
    q4=a34*b43;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c33=w1+w2+w3+w4;
    
    q1=a31*b14;
    q2=a32*b24;
    q3=a33*b34;
    q4=a34*b44;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c34=w1+w2+w3+w4;
    
    q1=a41*b11;
    q2=a42*b21;
    q3=a43*b31;
    q4=a44*b41;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c41=w1+w2+w3+w4;
    
    q1=a41*b12;
    q2=a42*b22;
    q3=a43*b32;
    q4=a44*b42;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c42=w1+w2+w3+w4;
    
    q1=a41*b13;
    q2=a42*b23;
    q3=a43*b33;
    q4=a44*b43;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c43=w1+w2+w3+w4;
    
    q1=a41*b14;
    q2=a42*b24;
    q3=a43*b34;
    q4=a44*b44;
    q5={{16{q1[47]}},q1[47:15]};
    w1=q5[23:0];
    q5={{16{q2[47]}},q2[47:15]};
    w2=q5[23:0];
    q5={{16{q3[47]}},q3[47:15]};
    w3=q5[23:0];
    q5={{16{q4[47]}},q4[47:15]};
    w4=q5[23:0];
    c44=w1+w2+w3+w4;

end
endmodule