module ml_22(

	input wire signed [23:0] a,b,c,d,a1,b1,c1,d1,

	output reg signed [23:0] b11,b12,b21,b22
);

reg signed [47:0] q1,q2,q3,q4;
reg signed [23:0] w1,w2;

always @(*) 
begin
    q1=a*a1;
    q2={{16{q1[47]}},q1[47:15]};
    w1=q2[23:0];
    q1=b*c1;
    q2={{16{q1[47]}},q1[47:15]};
    w2=q2[23:0];
    b11=w1+w2;
    
    q1=a*b1;
    q2={{16{q1[47]}},q1[47:15]};
    w1=q2[23:0];
    q1=b*d1;
    q2={{16{q1[47]}},q1[47:15]};
    w2=q2[23:0];
    b12=w1+w2;
    
    q1=c*a1;
    q2={{16{q1[47]}},q1[47:15]};
    w1=q2[23:0];
    q1=d*c1;
    q2={{16{q1[47]}},q1[47:15]};
    w2=q2[23:0];
    b21=w1+w2;
    
    q1=c*b1;
    q2={{16{q1[47]}},q1[47:15]};
    w1=q2[23:0];
    q1=d*d1;
    q2={{16{q1[47]}},q1[47:15]};
    w2=q2[23:0];
    b22=w1+w2;

end
endmodule
