// `include "../include/AXI_define.svh"

// `include "../../src/AXI/ReadControl.sv"
// `include "../../src/AXI/WriteControl.sv"

// `include "../../src/AXI/AFIFO/AFIFO_Rx.sv"
// `include "../../src/AXI/AFIFO/AFIFO_Tx.sv"
// `include "../../src/AXI/AFIFO/Vector_SYNC.sv"

module AXI(
input logic                       CPU_CLK_i,     
input logic                       AXI_CLK_i,        
input logic                       ROM_CLK_i,      
input logic                       DRAM_CLK_i,
input logic                       SRAM_CLK_i,
input logic                       DMA_CLK_i,
input logic                       WDT_CLK_i,
input logic                       CPU_RST_i,      
input logic                       AXI_RST_i,        
input logic                       ROM_RST_i,      
input logic                       DRAM_RST_i,
input logic                       SRAM_RST_i,           
input logic                       DMA_RST_i,  
input logic                       WDT_RST_i,                  
//MASTER INTERFACE
// M0
// READ
input  logic [`AXI_ID_BITS-1:0]   ARID_M0,
input  logic [`AXI_ADDR_BITS-1:0] ARADDR_M0,
input  logic [`AXI_LEN_BITS-1:0]  ARLEN_M0,
input  logic [`AXI_SIZE_BITS-1:0] ARSIZE_M0,
input  logic [1:0]                ARBURST_M0,
input  logic                      ARVALID_M0,
output logic                      ARREADY_M0,
output logic [`AXI_ID_BITS-1:0]   RID_M0,
output logic [`AXI_DATA_BITS-1:0] RDATA_M0,
output logic [1:0]                RRESP_M0,
output logic                      RLAST_M0,
output logic                      RVALID_M0,
input  logic                      RREADY_M0,
// M1
// WRITE
input  logic[`AXI_ID_BITS-1:0]    AWID_M1,
input  logic[`AXI_ADDR_BITS-1:0]  AWADDR_M1,
input  logic[`AXI_LEN_BITS-1:0]   AWLEN_M1,
input  logic[`AXI_SIZE_BITS-1:0]  AWSIZE_M1,
input  logic[1:0]                 AWBURST_M1,
input  logic                      AWVALID_M1,
output logic                      AWREADY_M1,
input  logic [`AXI_DATA_BITS-1:0] WDATA_M1,
input  logic [`AXI_STRB_BITS-1:0] WSTRB_M1,
input  logic                      WLAST_M1,
input  logic                      WVALID_M1,
output logic                      WREADY_M1,
output logic [`AXI_ID_BITS-1:0]   BID_M1,
output logic [1:0]                BRESP_M1,
output logic                      BVALID_M1,
input  logic                      BREADY_M1,
// READ
input  logic [`AXI_ID_BITS-1:0]   ARID_M1,
input  logic [`AXI_ADDR_BITS-1:0] ARADDR_M1,
input  logic [`AXI_LEN_BITS-1:0]  ARLEN_M1,
input  logic [`AXI_SIZE_BITS-1:0] ARSIZE_M1,
input  logic [1:0]                ARBURST_M1,
input  logic                      ARVALID_M1,
output logic                      ARREADY_M1,
output logic [`AXI_ID_BITS-1:0]   RID_M1,
output logic [`AXI_DATA_BITS-1:0] RDATA_M1,
output logic [1:0]                RRESP_M1,
output logic                      RLAST_M1,
output logic                      RVALID_M1,
input  logic                      RREADY_M1,
// M2
// WRITE
input  logic[`AXI_ID_BITS-1:0]    AWID_M2,
input  logic[`AXI_ADDR_BITS-1:0]  AWADDR_M2,
input  logic[`AXI_LEN_BITS-1:0]   AWLEN_M2,
input  logic[`AXI_SIZE_BITS-1:0]  AWSIZE_M2,
input  logic[1:0]                 AWBURST_M2,
input  logic                      AWVALID_M2,
output logic                      AWREADY_M2,
input  logic [`AXI_DATA_BITS-1:0] WDATA_M2,
input  logic [`AXI_STRB_BITS-1:0] WSTRB_M2,
input  logic                      WLAST_M2,
input  logic                      WVALID_M2,
output logic                      WREADY_M2,
output logic [`AXI_ID_BITS-1:0]   BID_M2,
output logic [1:0]                BRESP_M2,
output logic                      BVALID_M2,
input  logic                      BREADY_M2,
// READ
input  logic [`AXI_ID_BITS-1:0]   ARID_M2,
input  logic [`AXI_ADDR_BITS-1:0] ARADDR_M2,
input  logic [`AXI_LEN_BITS-1:0]  ARLEN_M2,
input  logic [`AXI_SIZE_BITS-1:0] ARSIZE_M2,
input  logic [1:0]                ARBURST_M2,
input  logic                      ARVALID_M2,
output logic                      ARREADY_M2,
output logic [`AXI_ID_BITS-1:0]   RID_M2,
output logic [`AXI_DATA_BITS-1:0] RDATA_M2,
output logic [1:0]                RRESP_M2,
output logic                      RLAST_M2,
output logic                      RVALID_M2,
input  logic                      RREADY_M2,
//SLAVE INTERFACE
// S0
// READ
output logic [`AXI_IDS_BITS-1:0]  ARID_S0,
output logic[`AXI_ADDR_BITS-1:0]  ARADDR_S0,
output logic[`AXI_LEN_BITS-1:0]   ARLEN_S0,
output logic[`AXI_SIZE_BITS-1:0]  ARSIZE_S0,
output logic[1:0]                 ARBURST_S0,
output logic                      ARVALID_S0,
input  logic                      ARREADY_S0,
input  logic[`AXI_IDS_BITS-1:0]   RID_S0,
input  logic[`AXI_DATA_BITS-1:0]  RDATA_S0,
input  logic[1:0]                 RRESP_S0,
input  logic                      RLAST_S0,
input  logic                      RVALID_S0,
output logic                      RREADY_S0,
// S1
// WRITE
output logic [`AXI_IDS_BITS-1:0]  AWID_S1,
output logic[`AXI_ADDR_BITS-1:0]  AWADDR_S1,
output logic[`AXI_LEN_BITS-1:0]   AWLEN_S1,
output logic[`AXI_SIZE_BITS-1:0]  AWSIZE_S1,
output logic[1:0]                 AWBURST_S1,
output logic                      AWVALID_S1,
input  logic                      AWREADY_S1,
output logic [`AXI_DATA_BITS-1:0] WDATA_S1,
output logic [`AXI_STRB_BITS-1:0] WSTRB_S1,
output logic                      WLAST_S1,
output logic                      WVALID_S1,
input  logic                      WREADY_S1,
input  logic[`AXI_IDS_BITS-1:0]   BID_S1,
input  logic[1:0]                 BRESP_S1,
input  logic                      BVALID_S1,
output logic                      BREADY_S1,
// READ
output logic [`AXI_IDS_BITS-1:0]  ARID_S1,
output logic[`AXI_ADDR_BITS-1:0]  ARADDR_S1,
output logic[`AXI_LEN_BITS-1:0]   ARLEN_S1,
output logic[`AXI_SIZE_BITS-1:0]  ARSIZE_S1,
output logic[1:0]                 ARBURST_S1,
output logic                      ARVALID_S1,
input  logic                      ARREADY_S1,
input  logic[`AXI_IDS_BITS-1:0]   RID_S1,
input  logic[`AXI_DATA_BITS-1:0]  RDATA_S1,
input  logic[1:0]                 RRESP_S1,
input  logic                      RLAST_S1,
input  logic                      RVALID_S1,
output logic                      RREADY_S1,
// S2
// WRITE
output logic [`AXI_IDS_BITS-1:0]  AWID_S2,
output logic[`AXI_ADDR_BITS-1:0]  AWADDR_S2,
output logic[`AXI_LEN_BITS-1:0]   AWLEN_S2,
output logic[`AXI_SIZE_BITS-1:0]  AWSIZE_S2,
output logic[1:0]                 AWBURST_S2,
output logic                      AWVALID_S2,
input  logic                      AWREADY_S2,
output logic [`AXI_DATA_BITS-1:0] WDATA_S2,
output logic [`AXI_STRB_BITS-1:0] WSTRB_S2,
output logic                      WLAST_S2,
output logic                      WVALID_S2,
input  logic                      WREADY_S2,
input  logic [`AXI_IDS_BITS-1:0]  BID_S2,
input  logic [1:0]                BRESP_S2,
input  logic                      BVALID_S2,
output logic                      BREADY_S2,
// READ
output logic [`AXI_IDS_BITS-1:0]  ARID_S2,
output logic[`AXI_ADDR_BITS-1:0]  ARADDR_S2,
output logic[`AXI_LEN_BITS-1:0]   ARLEN_S2,
output logic[`AXI_SIZE_BITS-1:0]  ARSIZE_S2,
output logic [1:0]                ARBURST_S2,
output logic                      ARVALID_S2,
input  logic                      ARREADY_S2,
input  logic[`AXI_IDS_BITS-1:0]   RID_S2,
input  logic[`AXI_DATA_BITS-1:0]  RDATA_S2,
input  logic[1:0]                 RRESP_S2,
input  logic                      RLAST_S2,
input  logic                      RVALID_S2,
output logic                      RREADY_S2,
// S3
// WRITE
output logic [`AXI_IDS_BITS-1:0]  AWID_S3,
output logic [`AXI_ADDR_BITS-1:0] AWADDR_S3,
output logic [`AXI_LEN_BITS-1:0]  AWLEN_S3,
output logic [`AXI_SIZE_BITS-1:0] AWSIZE_S3,
output logic [1:0]                AWBURST_S3,
output logic                      AWVALID_S3,
input  logic                      AWREADY_S3,
output logic [`AXI_DATA_BITS-1:0] WDATA_S3,
output logic [`AXI_STRB_BITS-1:0] WSTRB_S3,
output logic                      WLAST_S3,
output logic                      WVALID_S3,
input  logic                      WREADY_S3,
input  logic [`AXI_IDS_BITS-1:0]  BID_S3,
input  logic [1:0]                BRESP_S3,
input  logic                      BVALID_S3,
output logic                      BREADY_S3,
// READ
output logic [`AXI_IDS_BITS-1:0]  ARID_S3,
output logic [`AXI_ADDR_BITS-1:0] ARADDR_S3,
output logic [`AXI_LEN_BITS-1:0]  ARLEN_S3,
output logic [`AXI_SIZE_BITS-1:0] ARSIZE_S3,
output logic [1:0]                ARBURST_S3,
output logic                      ARVALID_S3,
input  logic                      ARREADY_S3,
input  logic [`AXI_IDS_BITS-1:0]  RID_S3,
input  logic [`AXI_DATA_BITS-1:0] RDATA_S3,
input  logic [1:0]                RRESP_S3,
input  logic                      RLAST_S3,
input  logic                      RVALID_S3,
output logic                      RREADY_S3,
// S4
// WRITE
output logic [`AXI_IDS_BITS-1:0]  AWID_S4,
output logic[`AXI_ADDR_BITS-1:0]  AWADDR_S4,
output logic[`AXI_LEN_BITS-1:0]   AWLEN_S4,
output logic[`AXI_SIZE_BITS-1:0]  AWSIZE_S4,
output logic[1:0]                 AWBURST_S4,
output logic                      AWVALID_S4,
input  logic                      AWREADY_S4,
output logic [`AXI_DATA_BITS-1:0] WDATA_S4,
output logic [`AXI_STRB_BITS-1:0] WSTRB_S4,
output logic                      WLAST_S4,
output logic                      WVALID_S4,
input  logic                      WREADY_S4,
input  logic[`AXI_IDS_BITS-1:0]   BID_S4,
input  logic[1:0]                 BRESP_S4,
input  logic                      BVALID_S4,
output logic                      BREADY_S4,
// READ
output logic [`AXI_IDS_BITS-1:0]  ARID_S4,
output logic[`AXI_ADDR_BITS-1:0]  ARADDR_S4,
output logic[`AXI_LEN_BITS-1:0]   ARLEN_S4,
output logic[`AXI_SIZE_BITS-1:0]  ARSIZE_S4,
output logic[1:0]                 ARBURST_S4,
output logic                      ARVALID_S4,
input  logic                      ARREADY_S4,
input  logic[`AXI_IDS_BITS-1:0]   RID_S4,
input  logic[`AXI_DATA_BITS-1:0]  RDATA_S4,
input  logic[1:0]                 RRESP_S4,
input  logic                      RLAST_S4,
input  logic                      RVALID_S4,
output logic                      RREADY_S4,
// S5
// WRITE
output logic [`AXI_IDS_BITS-1:0]  AWID_S5,
output logic [`AXI_ADDR_BITS-1:0] AWADDR_S5,
output logic [`AXI_LEN_BITS-1:0]  AWLEN_S5,
output logic [`AXI_SIZE_BITS-1:0] AWSIZE_S5,
output logic [1:0]                AWBURST_S5,
output logic                      AWVALID_S5,
input  logic                      AWREADY_S5,
output logic [`AXI_DATA_BITS-1:0] WDATA_S5,
output logic [`AXI_STRB_BITS-1:0] WSTRB_S5,
output logic                      WLAST_S5,
output logic                      WVALID_S5,
input  logic                      WREADY_S5,
input  logic [`AXI_IDS_BITS-1:0]  BID_S5,
input logic [1:0]                 BRESP_S5,
input logic                       BVALID_S5,
output logic                      BREADY_S5,
// READ
output logic [`AXI_IDS_BITS-1:0]  ARID_S5,
output logic [`AXI_ADDR_BITS-1:0] ARADDR_S5,
output logic [`AXI_LEN_BITS-1:0]  ARLEN_S5,
output logic [`AXI_SIZE_BITS-1:0] ARSIZE_S5,
output logic [1:0]                ARBURST_S5,
output logic                      ARVALID_S5,
input  logic                      ARREADY_S5,
input  logic [`AXI_IDS_BITS-1:0]  RID_S5,
input  logic [`AXI_DATA_BITS-1:0] RDATA_S5,
input  logic [1:0]                RRESP_S5,
input  logic                      RLAST_S5,
input  logic                      RVALID_S5,
output logic                      RREADY_S5
  
);



/////////////////////////////////////
	ReadControl read0
	(
		// .clk(AXI_CLK_i),
		// .rst(AXI_RST_i),
		.CPU_CLK_i 	(CPU_CLK_i ),
		.AXI_CLK_i 	(AXI_CLK_i ),
		.ROM_CLK_i 	(ROM_CLK_i ),
		.DRAM_CLK_i	(DRAM_CLK_i),
		.SRAM_CLK_i	(SRAM_CLK_i),
		.DMA_CLK_i	(DMA_CLK_i),
		.WDT_CLK_i	(WDT_CLK_i),
		.CPU_RST_i 	(CPU_RST_i ),
		.AXI_RST_i 	(AXI_RST_i ),
		.ROM_RST_i 	(ROM_RST_i ),
		.DRAM_RST_i	(DRAM_RST_i),
		.SRAM_RST_i	(SRAM_RST_i),
		.DMA_RST_i	(DMA_RST_i),
		.WDT_RST_i	(WDT_RST_i),
		// Master
		// READ ADDRESS0
		.ARID_M0(ARID_M0),
		.ARADDR_M0(ARADDR_M0),
		.ARLEN_M0(ARLEN_M0),
		.ARSIZE_M0(ARSIZE_M0),
		.ARBURST_M0(ARBURST_M0),
		.ARVALID_M0(ARVALID_M0),
		.ARREADY_M0(ARREADY_M0),
		// READ DATA0
		.RID_M0(RID_M0),
		.RDATA_M0(RDATA_M0),
		.RRESP_M0(RRESP_M0),
		.RLAST_M0(RLAST_M0),
		.RVALID_M0(RVALID_M0),
		.RREADY_M0(RREADY_M0),
		// READ ADDRESS1
		.ARID_M1(ARID_M1),
		.ARADDR_M1(ARADDR_M1),
		.ARLEN_M1(ARLEN_M1),
		.ARSIZE_M1(ARSIZE_M1),
		.ARBURST_M1(ARBURST_M1),
		.ARVALID_M1(ARVALID_M1),
		.ARREADY_M1(ARREADY_M1),
		// READ DATA1
		.RID_M1(RID_M1),
		.RDATA_M1(RDATA_M1),
		.RRESP_M1(RRESP_M1),
		.RLAST_M1(RLAST_M1),
		.RVALID_M1(RVALID_M1),
		.RREADY_M1(RREADY_M1),
		// READ ADDRESS2
		.ARID_M2(ARID_M2),
		.ARADDR_M2(ARADDR_M2),
		.ARLEN_M2(ARLEN_M2),
		.ARSIZE_M2(ARSIZE_M2),
		.ARBURST_M2(ARBURST_M2),
		.ARVALID_M2(ARVALID_M2),
		.ARREADY_M2(ARREADY_M2),
		// READ DATA2
		.RID_M2(RID_M2),
		.RDATA_M2(RDATA_M2),
		.RRESP_M2(RRESP_M2),
		.RLAST_M2(RLAST_M2),
		.RVALID_M2(RVALID_M2),
		.RREADY_M2(RREADY_M2),

		// Slave
		///// READ ADDRESS S0 (ROM)/////
		.ARID_S0(ARID_S0),
		.ARADDR_S0(ARADDR_S0),
		.ARLEN_S0(ARLEN_S0),
		.ARSIZE_S0(ARSIZE_S0),
		.ARBURST_S0(ARBURST_S0),
		.ARVALID_S0(ARVALID_S0),
		.ARREADY_S0(ARREADY_S0),
		// READ DATA S0
		.RID_S0(RID_S0),
		.RDATA_S0(RDATA_S0),
		.RRESP_S0(RRESP_S0),
		.RLAST_S0(RLAST_S0),
		.RVALID_S0(RVALID_S0),
		.RREADY_S0(RREADY_S0),
		///// READ ADDRESS S1 (IM SRAM)/////
		.ARID_S1(ARID_S1),
		.ARADDR_S1(ARADDR_S1),
		.ARLEN_S1(ARLEN_S1),
		.ARSIZE_S1(ARSIZE_S1),
		.ARBURST_S1(ARBURST_S1),
		.ARVALID_S1(ARVALID_S1),
		.ARREADY_S1(ARREADY_S1),
		// READ DATA S1
		.RID_S1(RID_S1),
		.RDATA_S1(RDATA_S1),
		.RRESP_S1(RRESP_S1),
		.RLAST_S1(RLAST_S1),
		.RVALID_S1(RVALID_S1),
		.RREADY_S1(RREADY_S1),
		///// READ ADDRESS S2 (DM SRAM)/////
		.ARID_S2(ARID_S2),
		.ARADDR_S2(ARADDR_S2),
		.ARLEN_S2(ARLEN_S2),
		.ARSIZE_S2(ARSIZE_S2),
		.ARBURST_S2(ARBURST_S2),
		.ARVALID_S2(ARVALID_S2),
		.ARREADY_S2(ARREADY_S2),
		// READ DATA S2
		.RID_S2(RID_S2),
		.RDATA_S2(RDATA_S2),
		.RRESP_S2(RRESP_S2),
		.RLAST_S2(RLAST_S2),
		.RVALID_S2(RVALID_S2),
		.RREADY_S2(RREADY_S2),
		///// READ ADDRESS S3 (DMA)/////
		.ARID_S3(ARID_S3),
		.ARADDR_S3(ARADDR_S3),
		.ARLEN_S3(ARLEN_S3),
		.ARSIZE_S3(ARSIZE_S3),
		.ARBURST_S3(ARBURST_S3),
		.ARVALID_S3(ARVALID_S3),
		.ARREADY_S3(ARREADY_S3),
		// READ DATA S3
		.RID_S3(RID_S3),
		.RDATA_S3(RDATA_S3),
		.RRESP_S3(RRESP_S3),
		.RLAST_S3(RLAST_S3),
		.RVALID_S3(RVALID_S3),
		.RREADY_S3(RREADY_S3),
		///// READ ADDRESS S4 (WDT)/////
		.ARID_S4(ARID_S4),
		.ARADDR_S4(ARADDR_S4),
		.ARLEN_S4(ARLEN_S4),
		.ARSIZE_S4(ARSIZE_S4),
		.ARBURST_S4(ARBURST_S4),
		.ARVALID_S4(ARVALID_S4),
		.ARREADY_S4(ARREADY_S4),
		// READ DATA S4
		.RID_S4(RID_S4),
		.RDATA_S4(RDATA_S4),
		.RRESP_S4(RRESP_S4),
		.RLAST_S4(RLAST_S4),
		.RVALID_S4(RVALID_S4),
		.RREADY_S4(RREADY_S4),
		///// READ ADDRESS S5 (DRAM)/////
		.ARID_S5(ARID_S5),
		.ARADDR_S5(ARADDR_S5),
		.ARLEN_S5(ARLEN_S5),
		.ARSIZE_S5(ARSIZE_S5),
		.ARBURST_S5(ARBURST_S5),
		.ARVALID_S5(ARVALID_S5),
		.ARREADY_S5(ARREADY_S5),
		// READ DATA S5
		.RID_S5(RID_S5),
		.RDATA_S5(RDATA_S5),
		.RRESP_S5(RRESP_S5),
		.RLAST_S5(RLAST_S5),
		.RVALID_S5(RVALID_S5),
		.RREADY_S5(RREADY_S5)								
	);
    
	WriteControl write0
	(
		// .clk(AXI_CLK_i),
		// .rst(AXI_RST_i),
		.CPU_CLK_i 	(CPU_CLK_i ),
		.AXI_CLK_i 	(AXI_CLK_i ),
		.ROM_CLK_i 	(ROM_CLK_i ),
		.DRAM_CLK_i	(DRAM_CLK_i),
		.SRAM_CLK_i	(SRAM_CLK_i),
		.DMA_CLK_i	(DMA_CLK_i),
		.WDT_CLK_i	(WDT_CLK_i),
		.CPU_RST_i 	(CPU_RST_i ),
		.AXI_RST_i 	(AXI_RST_i ),
		.ROM_RST_i 	(ROM_RST_i ),
		.DRAM_RST_i	(DRAM_RST_i),
		.SRAM_RST_i	(SRAM_RST_i),
		.DMA_RST_i	(DMA_RST_i),
		.WDT_RST_i	(WDT_RST_i),

		// Master
		// WRITE ADDRESS1
		.AWID_M1(AWID_M1),
		.AWADDR_M1(AWADDR_M1),
		.AWLEN_M1(AWLEN_M1),
		.AWSIZE_M1(AWSIZE_M1),
		.AWBURST_M1(AWBURST_M1),
		.AWVALID_M1(AWVALID_M1),
		.AWREADY_M1(AWREADY_M1),
		// WRITE DATA1
		.WDATA_M1(WDATA_M1),
		.WSTRB_M1(WSTRB_M1),
		.WLAST_M1(WLAST_M1),
		.WVALID_M1(WVALID_M1),
		.WREADY_M1(WREADY_M1),
		// WRITE RESPONSE1
		.BID_M1(BID_M1),
		.BRESP_M1(BRESP_M1),
		.BVALID_M1(BVALID_M1),
		.BREADY_M1(BREADY_M1),

		// WRITE ADDRESS2
		.AWID_M2(AWID_M2),
		.AWADDR_M2(AWADDR_M2),
		.AWLEN_M2(AWLEN_M2),
		.AWSIZE_M2(AWSIZE_M2),
		.AWBURST_M2(AWBURST_M2),
		.AWVALID_M2(AWVALID_M2),
		.AWREADY_M2(AWREADY_M2),
		// WRITE DATA2
		.WDATA_M2(WDATA_M2),
		.WSTRB_M2(WSTRB_M2),
		.WLAST_M2(WLAST_M2),
		.WVALID_M2(WVALID_M2),
		.WREADY_M2(WREADY_M2),
		// WRITE RESPONSE2
		.BID_M2(BID_M2),
		.BRESP_M2(BRESP_M2),
		.BVALID_M2(BVALID_M2),
		.BREADY_M2(BREADY_M2),

		// Slave
		////// WRITE ADDRESS S1
		.AWID_S1(AWID_S1),
		.AWADDR_S1(AWADDR_S1),
		.AWLEN_S1(AWLEN_S1),
		.AWSIZE_S1(AWSIZE_S1),
		.AWBURST_S1(AWBURST_S1),
		.AWVALID_S1(AWVALID_S1),
		.AWREADY_S1(AWREADY_S1),
		// WRITE DATA S1
		.WDATA_S1(WDATA_S1),
		.WSTRB_S1(WSTRB_S1),
		.WLAST_S1(WLAST_S1),
		.WVALID_S1(WVALID_S1),
		.WREADY_S1(WREADY_S1),
		// WRITE RESPONSE S1
		.BID_S1(BID_S1),
		.BRESP_S1(BRESP_S1),
		.BVALID_S1(BVALID_S1),
		.BREADY_S1(BREADY_S1),
		////// WRITE ADDRESS S2
		.AWID_S2(AWID_S2),
		.AWADDR_S2(AWADDR_S2),
		.AWLEN_S2(AWLEN_S2),
		.AWSIZE_S2(AWSIZE_S2),
		.AWBURST_S2(AWBURST_S2),
		.AWVALID_S2(AWVALID_S2),
		.AWREADY_S2(AWREADY_S2),
		// WRITE DATA S2
		.WDATA_S2(WDATA_S2),
		.WSTRB_S2(WSTRB_S2),
		.WLAST_S2(WLAST_S2),
		.WVALID_S2(WVALID_S2),
		.WREADY_S2(WREADY_S2),
		// WRITE RESPONSE S2
		.BID_S2(BID_S2),
		.BRESP_S2(BRESP_S2),
		.BVALID_S2(BVALID_S2),
		.BREADY_S2(BREADY_S2),
		// WRITE ADDRESS S3 
		.AWID_S3(AWID_S3),
		.AWADDR_S3(AWADDR_S3),
		.AWLEN_S3(AWLEN_S3),
		.AWSIZE_S3(AWSIZE_S3),
		.AWBURST_S3(AWBURST_S3),
		.AWVALID_S3(AWVALID_S3),
		.AWREADY_S3(AWREADY_S3),
		// WRITE DATA S3
		.WDATA_S3(WDATA_S3),
		.WSTRB_S3(WSTRB_S3),
		.WLAST_S3(WLAST_S3),
		.WVALID_S3(WVALID_S3),
		.WREADY_S3(WREADY_S3),
		// WRITE RESPONSE1 S3
		.BID_S3(BID_S3),
		.BRESP_S3(BRESP_S3),
		.BVALID_S3(BVALID_S3),
		.BREADY_S3(BREADY_S3),
		// WRITE ADDRESS S4 
		.AWID_S4(AWID_S4),
		.AWADDR_S4(AWADDR_S4),
		.AWLEN_S4(AWLEN_S4),
		.AWSIZE_S4(AWSIZE_S4),
		.AWBURST_S4(AWBURST_S4),
		.AWVALID_S4(AWVALID_S4),
		.AWREADY_S4(AWREADY_S4),
		// WRITE DATA S4
		.WDATA_S4(WDATA_S4),
		.WSTRB_S4(WSTRB_S4),
		.WLAST_S4(WLAST_S4),
		.WVALID_S4(WVALID_S4),
		.WREADY_S4(WREADY_S4),
		// WRITE RESPONSE S4
		.BID_S4(BID_S4),
		.BRESP_S4(BRESP_S4),
		.BVALID_S4(BVALID_S4),
		.BREADY_S4(BREADY_S4),
		// WRITE ADDRESS S5 
		.AWID_S5(AWID_S5),
		.AWADDR_S5(AWADDR_S5),
		.AWLEN_S5(AWLEN_S5),
		.AWSIZE_S5(AWSIZE_S5),
		.AWBURST_S5(AWBURST_S5),
		.AWVALID_S5(AWVALID_S5),
		.AWREADY_S5(AWREADY_S5),
		// WRITE DATA S5
		.WDATA_S5(WDATA_S5),
		.WSTRB_S5(WSTRB_S5),
		.WLAST_S5(WLAST_S5),
		.WVALID_S5(WVALID_S5),
		.WREADY_S5(WREADY_S5),
		// WRITE RESP S5
		.BID_S5(BID_S5),
		.BRESP_S5(BRESP_S5),
		.BVALID_S5(BVALID_S5),
		.BREADY_S5(BREADY_S5)
	);


endmodule
